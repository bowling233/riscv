module ALU (
  input [31:0]  A,
  input [31:0]  B,
  input [2:0]   ALU_operation,
  output[31:0]  res,
  output        zero
);
// Your code

endmodule