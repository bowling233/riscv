`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/02/21 10:08:22
// Design Name: 
// Module Name: div32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module divider(
    input   clk,
    input   rst,
    input   start,
    input[31:0] dividend, 
    input[31:0] divisor,
    output divide_zero,
    output  finish,
    output[31:0] res,
    output[31:0] rem
); 
		
    
    
	endmodule

